LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY LOCKIS IS
PORT(le:IN STD_LOGIC;
		dd:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		qq:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END LOCKIS;
ARCHITECTURE one OF LOCKIS IS
BEGIN
	PROCESS (le,dd)
		BEGIN
			IF (le='1')THEN
				qq<=dd;
			END IF;
		END PROCESS;
	END one;